module or_ga(g_if inf);
  
  assign inf.dut.y=inf.dut.a|inf.dut.b;
  
endmodule
