class trans;
  bit clk;
  bit rst;
  randc bit D;
  bit Q;
endclass
